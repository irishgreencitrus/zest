module main

fn main() {
    println("HelloWorld!!")
}
